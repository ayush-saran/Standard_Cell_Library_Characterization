* SKY130 Spice File.

.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice"

.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice"

.include "../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"

.include "corners/tt/rf.spice"
.include "all.spice"
.include "corners/tt/nonfet.spice"

